module xor_memory(clk);
  input clk;

endmodule
